asczcasdasdsadsadasdsafsadfs