asczcasdasdsadsadasdsafsadfssadsada